library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;

library UNISIM;
use UNISIM.VComponents.ALL;

entity ROM_1024x16_DUO is
	port (
		-- CLOCK
		I_CLK	: in	STD_LOGIC;
		
		-- RESET
		I_RST	: in	STD_LOGIC;
		
		-- ADDRESS
		I_ADDR	: in	STD_LOGIC_VECTOR (9 downto 0);
		
		-- DUAL CHANNEL DATA
		O_DATA0	: out	STD_LOGIC_VECTOR (15 downto 0);
		O_DATA1	: out	STD_LOGIC_VECTOR (15 downto 0));
end ROM_1024x16_DUO;

architecture arch of ROM_1024x16_DUO is

	component ROM_512x16 is
		generic (	
		
			-- MEMORY MAP
			INIT_00	: BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_01	: BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_02	: BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_03	: BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_04	: BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_05	: BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_06	: BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_07	: BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_08	: BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_09	: BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_0A	: BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_0B	: BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_0C	: BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_0D	: BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_0E	: BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_0F	: BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_10	: BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_11	: BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_12	: BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_13	: BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_14	: BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_15	: BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_16	: BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_17	: BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_18	: BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_19	: BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_1A	: BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_1B	: BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_1C	: BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_1D	: BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_1E	: BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_1F	: BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000");
			
		port (
			-- CLOCK
			I_CLK	: in	STD_LOGIC;
			
			-- RESET
			I_RST	: in	STD_LOGIC;
			
			-- ADDRESS
			I_ADDR	: in	STD_LOGIC_VECTOR (8 downto 0);
			
			-- DATA
			O_DATA	: out	STD_LOGIC_VECTOR (15 downto 0));
	end component;	
	
	constant L_GND : STD_LOGIC := '0';
	
	type SLV2x16 is 
		array(0 to 1) of STD_LOGIC_VECTOR(15 downto 0);
	type SLV2x10 is 
		array(0 to 1) of STD_LOGIC_VECTOR(8 downto 0);
	
	signal ROM_out	: SLV2x16 := (others => (others => L_GND));
	signal ROM_addr	: SLV2x10 := (others => (others => L_GND));
	
	type SLV32x256 is 
		array(0 to 31) of bit_vector(255 downto 0);
	
	type SLV32x256_duo is 
		array(0 to 1) of SLV32x256;
		
	constant ROM_init : SLV32x256_duo := (
	
	(0 => X"0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0009_0007_0005_0003_0001",		
		others => X"0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000"),
			
	(0 => X"0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_000A_0008_0006_0004_0002",		
		others => X"0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000"));
		
	signal L_CLK : STD_LOGIC := '0';
begin

	process(I_CLK, I_ADDR)
		variable v_ROM_addr0 : STD_LOGIC_VECTOR(8 downto 0);
	begin
	
		if (I_ADDR(0)='0') then
			ROM_addr(0) <= I_ADDR(9 downto 1);
		else
			ROM_addr(0) <= conv_std_logic_vector(UNSIGNED(I_ADDR(9 downto 1))+1, ROM_addr(0)'length);
		end if;
		
		ROM_addr(1) <= I_ADDR(9 downto 1);
		
		L_CLK <= I_CLK;
	end process;
	
	MAIN : for i in 0 to 1
	generate
		ROM_UNIT: ROM_512x16
			generic map(
				INIT_00 => ROM_init(i)(0),
				INIT_01 => ROM_init(i)(1),
				INIT_02 => ROM_init(i)(2),
				INIT_03 => ROM_init(i)(3),
				INIT_04 => ROM_init(i)(4),
				INIT_05 => ROM_init(i)(5),
				INIT_06 => ROM_init(i)(6),
				INIT_07 => ROM_init(i)(7),
				INIT_08 => ROM_init(i)(8),
				INIT_09 => ROM_init(i)(9),
				INIT_0A => ROM_init(i)(10),
				INIT_0B => ROM_init(i)(11),
				INIT_0C => ROM_init(i)(12),
				INIT_0D => ROM_init(i)(13),
				INIT_0E => ROM_init(i)(14),
				INIT_0F => ROM_init(i)(15),
				INIT_10 => ROM_init(i)(16),
				INIT_11 => ROM_init(i)(17),
				INIT_12 => ROM_init(i)(18),
				INIT_13 => ROM_init(i)(19),
				INIT_14 => ROM_init(i)(20),
				INIT_15 => ROM_init(i)(21),
				INIT_16 => ROM_init(i)(22),
				INIT_17 => ROM_init(i)(23),
				INIT_18 => ROM_init(i)(24),
				INIT_19 => ROM_init(i)(25),
				INIT_1A => ROM_init(i)(26),
				INIT_1B => ROM_init(i)(27),
				INIT_1C => ROM_init(i)(28),
				INIT_1D => ROM_init(i)(29),
				INIT_1E => ROM_init(i)(30),
				INIT_1F => ROM_init(i)(31))				
			port map( 
				I_CLK 	=> L_CLK,
				I_RST 	=> I_RST,
				I_ADDR 	=> ROM_addr(i),
				O_DATA 	=> ROM_out(i));
	end generate;	
	
	OUTPUT : for i in 0 to 15
	generate
		MUX_OUT0: O_DATA0(i) <= ROM_out(
			conv_integer(
				NOT I_ADDR(0)))(i);
				
		MUX_OUT1: O_DATA1(i) <= ROM_out(
			conv_integer(
				I_ADDR(0)))(i);				
	end generate;
end arch;

