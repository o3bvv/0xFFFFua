library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;

library UNISIM;
use UNISIM.VComponents.ALL;

entity ROM_512x16 is
	generic (	
	
		-- MEMORY MAP
		INIT_00	: BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_01	: BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_02	: BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_03	: BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_04	: BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_05	: BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_06	: BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_07	: BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_08	: BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_09	: BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_0A	: BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_0B	: BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_0C	: BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_0D	: BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_0E	: BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_0F	: BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_10	: BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_11	: BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_12	: BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_13	: BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_14	: BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_15	: BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_16	: BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_17	: BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_18	: BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_19	: BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_1A	: BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_1B	: BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_1C	: BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_1D	: BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_1E	: BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_1F	: BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000");
		
	port (
		-- CLOCK
		I_CLK	: in	STD_LOGIC;
		
		-- RESET
		I_RST	: in	STD_LOGIC;
		
		-- ADDRESS
		I_ADDR	: in	STD_LOGIC_VECTOR (8 downto 0);
		
		-- DATA
		O_DATA	: out	STD_LOGIC_VECTOR (15 downto 0));
end ROM_512x16;

architecture arch of ROM_512x16 is

	component RAMB4_S16 is	
		generic (
			INIT_00 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_01 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_02 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_03 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_04 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_05 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_06 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_07 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_08 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_09 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_0A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_0B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_0C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_0D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_0E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_0F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000");
			
		port (
			DI	 : in  STD_LOGIC_VECTOR (15 downto 0);
			EN 	 : in  STD_ULOGIC;
			WE 	 : in  STD_ULOGIC;
			RST  : in  STD_ULOGIC;
			CLK  : in  STD_ULOGIC;
			ADDR : in  STD_LOGIC_VECTOR (7 downto 0);
			DO 	 : out STD_LOGIC_VECTOR (15 downto 0));
	end component;
	
	constant L_GND		: STD_LOGIC := '0';
	constant L_VCC		: STD_LOGIC := '1';
	constant L_GND_16	: STD_LOGIC_VECTOR(15 downto 0) := (others => L_GND);	
	
	type SLV2x16 is 
		array(0 to 1) of STD_LOGIC_VECTOR(15 downto 0);
	
	signal ROM_out	: SLV2x16 := (others => (others => L_GND));
	
	type SLV32x256 is 
		array(0 to 31) of bit_vector(255 downto 0);
	
	constant ROM_init : SLV32x256 := (
		INIT_00, INIT_01, INIT_02, INIT_03, INIT_04, INIT_05, INIT_07, INIT_07,
		INIT_08, INIT_09, INIT_0A, INIT_0B, INIT_0C, INIT_0D, INIT_0E, INIT_0F,
		INIT_10, INIT_11, INIT_12, INIT_13, INIT_14, INIT_15, INIT_17, INIT_17,
		INIT_18, INIT_19, INIT_1A, INIT_1B, INIT_1C, INIT_1D, INIT_1E, INIT_1F);
begin

	MAIN : for i in 0 to 1
	generate
		ROM_UNIT: RAMB4_S16 
			generic map(
				INIT_00 => ROM_init(16*i+0),
				INIT_01 => ROM_init(16*i+1),
				INIT_02 => ROM_init(16*i+2),
				INIT_03 => ROM_init(16*i+3),
				INIT_04 => ROM_init(16*i+4),
				INIT_05 => ROM_init(16*i+5),
				INIT_06 => ROM_init(16*i+6),
				INIT_07 => ROM_init(16*i+7),
				INIT_08 => ROM_init(16*i+8),
				INIT_09 => ROM_init(16*i+9),
				INIT_0A => ROM_init(16*i+10),
				INIT_0B => ROM_init(16*i+11),
				INIT_0C => ROM_init(16*i+12),
				INIT_0D => ROM_init(16*i+13),
				INIT_0E => ROM_init(16*i+14),
				INIT_0F => ROM_init(16*i+15))
			port map (
				CLK		=> I_CLK,
				RST 	=> I_RST,
				EN		=> L_VCC,
				WE 		=> L_GND,
				DI		=> L_GND_16,
				ADDR 	=> I_ADDR(7 downto 0),
				DO 		=> ROM_out(i));
	end generate;

	OUTPUT : for i in 0 to 15 generate
		MUX_OUT: O_DATA(i) <= ROM_out(
			conv_integer(
				I_ADDR(8)))(i);
	end generate;
end arch;

