--------------------------------------------------------------------------------
-- Instructions ROM
-- 1Kx16bit
--------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

library UNISIM;
use UNISIM.VComponents.all;

entity ROM1Kx16 is
	generic (
		INIT_00	: bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_01	: bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_02	: bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_03	: bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_04	: bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_05	: bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_06	: bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_07	: bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_08	: bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_09	: bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_0A	: bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_0B	: bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_0C	: bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_0D	: bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_0E	: bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_0F	: bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_10	: bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_11	: bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_12	: bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_13	: bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_14	: bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_15	: bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_16	: bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_17	: bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_18	: bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_19	: bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_1A	: bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_1B	: bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_1C	: bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_1D	: bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_1E	: bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_1F	: bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_20	: bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_21	: bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_22	: bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_23	: bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_24	: bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_25	: bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_26	: bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_27	: bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_28	: bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_29	: bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_2A	: bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_2B	: bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_2C	: bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_2D	: bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_2E	: bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_2F	: bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_30	: bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_31	: bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_32	: bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_33	: bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_34	: bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_35	: bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_36	: bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_37	: bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_38	: bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_39	: bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_3A	: bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_3B	: bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_3C	: bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_3D	: bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_3E	: bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
		INIT_3F	: bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000");
	port ( 
		I_CLK 	: in	STD_LOGIC;
		I_RST 	: in	STD_LOGIC;
		I_ADDR 	: in	STD_LOGIC_VECTOR (9 downto 0);
		O_DATA 	: out	STD_LOGIC_VECTOR (15 downto 0));
end ROM1Kx16;

architecture struct of ROM1Kx16 is
	
	component MUX4 is
		port ( 
			I0 		: in  STD_LOGIC;
			I1 		: in  STD_LOGIC;
			I2 		: in  STD_LOGIC;
			I3 		: in  STD_LOGIC;
			I_ADDR 	: in  STD_LOGIC_VECTOR (1 downto 0);
			O		: out STD_LOGIC);
	end component;
		
	component RAMB4_S16 is
	
		generic (
			INIT_00 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_01 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_02 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_03 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_04 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_05 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_06 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_07 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_08 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_09 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_0A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_0B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_0C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_0D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_0E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
			INIT_0F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000");
			
		port (
			DI: in STD_LOGIC_VECTOR (15 downto 0);
			EN : in STD_ULOGIC;
			WE : in STD_ULOGIC;
			RST : in STD_ULOGIC;
			CLK : in STD_ULOGIC;
			ADDR: in STD_LOGIC_VECTOR (7 downto 0);
			DO : out STD_LOGIC_VECTOR (15 downto 0));
	end component;
	
	type SLV4x16 is 
		array(0 to 3) of STD_LOGIC_VECTOR(15 downto 0);
	
	signal ROM_out	: SLV4x16;	

	constant L_GND_16	: STD_LOGIC_VECTOR(15 downto 0) := (others => '0');
	constant L_GND		: STD_LOGIC := '0';
	constant L_VCC		: STD_LOGIC := '1';
	
	type SLV64x256 is 
		array(0 to 63) of bit_vector(255 downto 0);
	
	constant ROM_init : SLV64x256 := (
		INIT_00, INIT_01, INIT_02, INIT_03, INIT_04, INIT_05, INIT_07, INIT_07,
		INIT_08, INIT_09, INIT_0A, INIT_0B, INIT_0C, INIT_0D, INIT_0E, INIT_0F,
		INIT_10, INIT_11, INIT_12, INIT_13, INIT_14, INIT_15, INIT_17, INIT_17,
		INIT_18, INIT_19, INIT_1A, INIT_1B, INIT_1C, INIT_1D, INIT_1E, INIT_1F,
		INIT_20, INIT_21, INIT_22, INIT_23, INIT_24, INIT_25, INIT_27, INIT_27,
		INIT_28, INIT_29, INIT_2A, INIT_2B, INIT_2C, INIT_2D, INIT_2E, INIT_2F,
		INIT_30, INIT_31, INIT_32, INIT_33, INIT_34, INIT_35, INIT_37, INIT_37,
		INIT_38, INIT_39, INIT_3A, INIT_3B, INIT_3C, INIT_3D, INIT_3E, INIT_3F);
begin
		
	MAIN : for i in 0 to 3
	generate
		ROM_UNIT: RAMB4_S16 
			generic map(
				INIT_00 => ROM_init(16*i+0),
				INIT_01 => ROM_init(16*i+1),
				INIT_02 => ROM_init(16*i+2),
				INIT_03 => ROM_init(16*i+3),
				INIT_04 => ROM_init(16*i+4),
				INIT_05 => ROM_init(16*i+5),
				INIT_06 => ROM_init(16*i+6),
				INIT_07 => ROM_init(16*i+7),
				INIT_08 => ROM_init(16*i+8),
				INIT_09 => ROM_init(16*i+9),
				INIT_0A => ROM_init(16*i+10),
				INIT_0B => ROM_init(16*i+11),
				INIT_0C => ROM_init(16*i+12),
				INIT_0D => ROM_init(16*i+13),
				INIT_0E => ROM_init(16*i+14),
				INIT_0F => ROM_init(16*i+15))
			port map (
				CLK		=> I_CLK,
				RST 	=> I_RST,
				EN		=> L_VCC,
				WE 		=> L_GND,
				DI		=> L_GND_16,
				ADDR 	=> I_ADDR(7 downto 0),
				DO 		=> ROM_out(i));
	end generate;
		
	OUTPUT : for i in 0 to 15 generate
		MUX_UNIT: MUX4
			port map (
				I3		=> ROM_out(3)(i),
				I2		=> ROM_out(2)(i),
				I1		=> ROM_out(1)(i),
				I0		=> ROM_out(0)(i),
				I_ADDR	=> I_ADDR(9 downto 8),
				O 		=> O_DATA(i));
	end generate;
end struct;

